package ieee_1149_tb_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ieee_1149_10_seq_item.sv"
`include "ieee_1149_10_sequence_lib.sv"
`include "ieee_1149_10_sequencer.sv"
`include "ieee_1149_10_driver.sv"
`include "ieee_1149_10_monitor.sv"
`include "ieee_1149_10_agent.sv"
`include "ieee_1149_10_virtual_sequencer.sv"
//`include "ieee_1149_10_coverage.sv"
`include "ieee_1149_10_scoreboard.sv"
`include "ieee_1149_10_env.sv"
`include "ieee_1149_10_virtual_sequence.sv"
`include "ieee_1149_10_test_lib.sv"
endpackage:ieee_1149_tb_pkg
